`include "sysconfig.v"
// 32位 Booth 华莱士乘法树，采用全加器（CSA）实现
module alu_mul_wallace_csa_32 (
    input                            clk,
    input                            rst,
    input                            rs1_signed_valid_i,
    input                            rs2_signed_valid_i,
    input  [  `XLEN_BUS] rs1_data_i,  // 32位
    input  [  `XLEN_BUS] rs2_data_i,  // 32位
    input                            mul_valid_i,
    output                           mul_ready_o,
    output [63:0]                    mul_out_o    // 64位输出
);

  // 寄存器已经复位
  localparam STATE_LEN = 3;
  localparam MUL_RST = 3'd0;
  localparam MUL_IDLE = 3'd1;
  localparam MUL_WAIT = 3'd3;

  wire _mul_valid = mul_valid_i;
  reg [STATE_LEN-1:0] mul_state;

  reg [2:0] mul_count;  // 减少计数位宽
  wire [2:0] mul_count_plus1 = mul_count + 'd1;

  reg mul_ready;
  reg [63:0] mul_data64;  // 64位结果

  reg [`XLEN_BUS] booth_rs1;
  reg [`XLEN_BUS] booth_rs2;
  reg booth_rs1_signed_valid;
  reg booth_rs2_signed_valid;

  wire [63:0] mul_final64;
  assign mul_ready_o = mul_ready;
  assign mul_out_o   = mul_data64;

  /* 乘法状态机切换 */
  always @(posedge clk) begin
    if (rst) begin
      mul_state <= MUL_RST;
      mul_ready <= `FALSE;
      mul_data64 <= 'b0;
      mul_count <= 'b0;
      booth_rs1 <= 'b0;
      booth_rs2 <= 'b0;
      booth_rs1_signed_valid <= 'b0;
      booth_rs2_signed_valid <= 'b0;
    end else begin
      case (mul_state)
        MUL_RST: begin
          mul_state <= MUL_IDLE;
        end
        MUL_IDLE: begin
          mul_ready <= `FALSE;
          mul_count <= 'b0;
          if (_mul_valid) begin  // 乘法请求
            mul_state <= MUL_WAIT;
            booth_rs1 <= rs1_data_i;
            booth_rs2 <= rs2_data_i;
            booth_rs1_signed_valid <= rs1_signed_valid_i;
            booth_rs2_signed_valid <= rs2_signed_valid_i;
          end
        end
        MUL_WAIT: begin
          if (~_mul_valid) begin
            mul_state <= MUL_IDLE;
          end else begin
            mul_count <= mul_count_plus1;
            if (mul_count == 'd2) begin  // 减少等待周期
              mul_data64 <= mul_final64;
              mul_state   <= MUL_IDLE;
              mul_ready   <= `TRUE;
            end
          end
        end
        default: begin
        end
      endcase
    end
  end

  wire [63:0] Partial_product[17-1:0];  // 32位需要17个部分积
  alu_mul_booth_r4_32 u_alu_mul_booth_r4_32 (
      .rs1_signed_valid_i(booth_rs1_signed_valid),
      .rs2_signed_valid_i(booth_rs2_signed_valid),
      .rs1_data_i        (booth_rs1),
      .rs2_data_i        (booth_rs2),
      .pp0_o             (Partial_product[0]),
      .pp1_o             (Partial_product[1]),
      .pp2_o             (Partial_product[2]),
      .pp3_o             (Partial_product[3]),
      .pp4_o             (Partial_product[4]),
      .pp5_o             (Partial_product[5]),
      .pp6_o             (Partial_product[6]),
      .pp7_o             (Partial_product[7]),
      .pp8_o             (Partial_product[8]),
      .pp9_o             (Partial_product[9]),
      .pp10_o            (Partial_product[10]),
      .pp11_o            (Partial_product[11]),
      .pp12_o            (Partial_product[12]),
      .pp13_o            (Partial_product[13]),
      .pp14_o            (Partial_product[14]),
      .pp15_o            (Partial_product[15]),
      .pp16_o            (Partial_product[16])
  );

  // 部分积生成 (共17个),缓存一个周期
  wire [63:0] step1_pp_q[17-1:0];

  genvar step1_Dflap;
  generate
    for (step1_Dflap = 0; step1_Dflap < 17; step1_Dflap = step1_Dflap + 1) begin
      regTemplate #(
          .WIDTH    (64),
          .RESET_VAL(0)
      ) u_regTemplate (
          .clk (clk),
          .rst (rst),
          .din (Partial_product[step1_Dflap]),
          .dout(step1_pp_q[step1_Dflap]),
          .wen (1'b1)
      );
    end
  endgenerate

  // 华莱士树压缩 - 32位版本需要更少的级数
  // 第一级: 17个部分积 -> 5个CSA(3-2) + 2个保留 = 12个输出
  localparam STEP1_CSA_NUM = 5;
  genvar step1_num_count;
  genvar step1_bit_count;
  wire [63:0] step1_sum  [STEP1_CSA_NUM-1:0];
  wire [63:0] step1_carry[STEP1_CSA_NUM-1:0];

  generate
    for (
        step1_num_count = 0; step1_num_count < STEP1_CSA_NUM; step1_num_count = step1_num_count + 1
    ) begin
      for (step1_bit_count = 0; step1_bit_count < 64; step1_bit_count = step1_bit_count + 1) begin
        full_adder u_full_adder_step1 (
            .a (step1_pp_q[step1_num_count*3+0][step1_bit_count]),
            .b (step1_pp_q[step1_num_count*3+1][step1_bit_count]),
            .ci(step1_pp_q[step1_num_count*3+2][step1_bit_count]),
            .s (step1_sum[step1_num_count][step1_bit_count]),
            .co(step1_carry[step1_num_count][step1_bit_count])
        );
      end
    end
  endgenerate

  // 第二级: 12个部分积 (5个和 + 5个进位 + 2个保留)
  wire [63:0] step2_pp_q[12-1:0];
  assign step2_pp_q[10] = step1_pp_q[15]; // 保留的两个部分积
  assign step2_pp_q[11] = step1_pp_q[16];
  
  genvar step2_pp_q_count;
  generate
    for (
        step2_pp_q_count = 0;
        step2_pp_q_count < STEP1_CSA_NUM;
        step2_pp_q_count = step2_pp_q_count + 1
    ) begin
      assign step2_pp_q[step2_pp_q_count*2+0] = step1_sum[step2_pp_q_count];
      assign step2_pp_q[step2_pp_q_count*2+1] = {step1_carry[step2_pp_q_count][62:0], 1'b0};
    end
  endgenerate

  // 第三级: 12个部分积 -> 4个CSA(3-2) = 8个输出
  localparam STEP2_CSA_NUM = 4;
  genvar step2_num_count;
  genvar step2_bit_count;
  wire [63:0] step2_sum  [STEP2_CSA_NUM-1:0];
  wire [63:0] step2_carry[STEP2_CSA_NUM-1:0];
  
  generate
    for (
        step2_num_count = 0; step2_num_count < STEP2_CSA_NUM; step2_num_count = step2_num_count + 1
    ) begin
      for (step2_bit_count = 0; step2_bit_count < 64; step2_bit_count = step2_bit_count + 1) begin
        full_adder u_full_adder_step2 (
            .a (step2_pp_q[step2_num_count*3+0][step2_bit_count]),
            .b (step2_pp_q[step2_num_count*3+1][step2_bit_count]),
            .ci(step2_pp_q[step2_num_count*3+2][step2_bit_count]),
            .s (step2_sum[step2_num_count][step2_bit_count]),
            .co(step2_carry[step2_num_count][step2_bit_count])
        );
      end
    end
  endgenerate

  // 第四级: 8个部分积 (4个和 + 4个进位)
  wire [63:0] step3_pp_q[8-1:0];
  genvar step3_pp_q_count;
  generate
    for (
        step3_pp_q_count = 0;
        step3_pp_q_count < STEP2_CSA_NUM;
        step3_pp_q_count = step3_pp_q_count + 1
    ) begin
      assign step3_pp_q[step3_pp_q_count*2+0] = step2_sum[step3_pp_q_count];
      assign step3_pp_q[step3_pp_q_count*2+1] = {step2_carry[step3_pp_q_count][62:0], 1'b0};
    end
  endgenerate

  // 第五级: 8个部分积 -> 2个CSA(3-2) + 2个保留 = 6个输出
  localparam STEP3_CSA_NUM = 2;
  genvar step3_num_count;
  genvar step3_bit_count;
  wire [63:0] step3_sum  [STEP3_CSA_NUM-1:0];
  wire [63:0] step3_carry[STEP3_CSA_NUM-1:0];
  
  generate
    for (
        step3_num_count = 0; step3_num_count < STEP3_CSA_NUM; step3_num_count = step3_num_count + 1
    ) begin
      for (step3_bit_count = 0; step3_bit_count < 64; step3_bit_count = step3_bit_count + 1) begin
        full_adder u_full_adder_step3 (
            .a (step3_pp_q[step3_num_count*3+0][step3_bit_count]),
            .b (step3_pp_q[step3_num_count*3+1][step3_bit_count]),
            .ci(step3_pp_q[step3_num_count*3+2][step3_bit_count]),
            .s (step3_sum[step3_num_count][step3_bit_count]),
            .co(step3_carry[step3_num_count][step3_bit_count])
        );
      end
    end
  endgenerate

  // 第六级: 6个部分积 (2个和 + 2个进位 + 2个保留)
  wire [63:0] step4_pp_q[6-1:0];
  assign step4_pp_q[4] = step3_pp_q[6]; // 保留的两个部分积
  assign step4_pp_q[5] = step3_pp_q[7];
  
  genvar step4_pp_q_count;
  generate
    for (
        step4_pp_q_count = 0;
        step4_pp_q_count < STEP3_CSA_NUM;
        step4_pp_q_count = step4_pp_q_count + 1
    ) begin
      assign step4_pp_q[step4_pp_q_count*2+0] = step3_sum[step4_pp_q_count];
      assign step4_pp_q[step4_pp_q_count*2+1] = {step3_carry[step4_pp_q_count][62:0], 1'b0};
    end
  endgenerate

  // 第七级: 6个部分积 -> 2个CSA(3-2) = 4个输出
  localparam STEP4_CSA_NUM = 2;
  genvar step4_num_count;
  genvar step4_bit_count;
  wire [63:0] step4_sum  [STEP4_CSA_NUM-1:0];
  wire [63:0] step4_carry[STEP4_CSA_NUM-1:0];
  
  generate
    for (
        step4_num_count = 0; step4_num_count < STEP4_CSA_NUM; step4_num_count = step4_num_count + 1
    ) begin
      for (step4_bit_count = 0; step4_bit_count < 64; step4_bit_count = step4_bit_count + 1) begin
        full_adder u_full_adder_step4 (
            .a (step4_pp_q[step4_num_count*3+0][step4_bit_count]),
            .b (step4_pp_q[step4_num_count*3+1][step4_bit_count]),
            .ci(step4_pp_q[step4_num_count*3+2][step4_bit_count]),
            .s (step4_sum[step4_num_count][step4_bit_count]),
            .co(step4_carry[step4_num_count][step4_bit_count])
        );
      end
    end
  endgenerate

  // 第八级: 4个部分积 -> 1个CSA(3-2) + 1个保留 = 3个输出
  wire [63:0] step5_pp_q[3-1:0];
  assign step5_pp_q[2] = step4_pp_q[5]; // 保留的部分积
  
  genvar step5_pp_q_count;
  generate
    for (
        step5_pp_q_count = 0;
        step5_pp_q_count < 1; // 只处理前两个
        step5_pp_q_count = step5_pp_q_count + 1
    ) begin
      assign step5_pp_q[step5_pp_q_count*2+0] = step4_sum[step5_pp_q_count];
      assign step5_pp_q[step5_pp_q_count*2+1] = {step4_carry[step5_pp_q_count][62:0], 1'b0};
    end
  endgenerate

  // 第九级: 3个部分积 -> 1个CSA(3-2) = 2个输出
  wire [63:0] step6_sum;
  wire [63:0] step6_carry;
  
  genvar step6_bit_count;
  generate
    for (step6_bit_count = 0; step6_bit_count < 64; step6_bit_count = step6_bit_count + 1) begin
      full_adder u_full_adder_step6 (
          .a (step5_pp_q[0][step6_bit_count]),
          .b (step5_pp_q[1][step6_bit_count]),
          .ci(step5_pp_q[2][step6_bit_count]),
          .s (step6_sum[step6_bit_count]),
          .co(step6_carry[step6_bit_count])
      );
    end
  endgenerate

  // 最终加法
  wire [63:0] step7_pp_a = step6_sum;
  wire [63:0] step7_pp_b = {step6_carry[62:0], 1'b0};
  
  // 插入流水线缓存
  wire [63:0] mul_final_a;
  wire [63:0] mul_final_b;
  regTemplate #(
      .WIDTH    (64),
      .RESET_VAL('b0)
  ) u_regTemplate_step7_a (
      .clk (clk),
      .rst (rst),
      .din (step7_pp_a),
      .dout(mul_final_a),
      .wen (1'b1)
  );
  regTemplate #(
      .WIDTH    (64),
      .RESET_VAL('b0)
  ) u_regTemplate_step7_b (
      .clk (clk),
      .rst (rst),
      .din (step7_pp_b),
      .dout(mul_final_b),
      .wen (1'b1)
  );

  /* 最终加法 */
  assign mul_final64 = mul_final_a + mul_final_b;

endmodule